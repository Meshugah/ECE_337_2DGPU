//Module: Request Unit
//Author(s): Noah Petersen
//Version: 1.0 Initial Design

module requestunit
(
	input wire primsel, //Will not need to use buffer for circle data
	input wire [31:0]buffdata, //Data from skeleton buffer, can be used as 
	input wire address,
	input wire dataready,
	output wire [4:0]sub_address,


);
/*
Requirements
	


*/


endmodule
