// $Id: $
// File name:   flex_stp_sr.sv
// Created:     9/13/2016
// Author:      Ahmad dit Ziad Dannawi
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: Flex serial to parallel shift register.
module flex_stp_sr
#(
 parameter NUM_BITS = 4,
 parameter SHIFT_MSB = 1
) 
(
 input wire clk, n_rst, shift_enable, serial_in,
 output wire [NUM_BITS-1:0]parallel_out
 ); 
   reg [NUM_BITS-1:0] 	temp_out;   
   genvar 			    i;

   always_ff @ (posedge clk, negedge n_rst)
     begin
	if (n_rst == 0) begin
	   temp_out <= {NUM_BITS{1'b1}};	   
	end else begin
	   if (shift_enable) begin
	      if (SHIFT_MSB) begin
	      	temp_out <= {temp_out[NUM_BITS-2:0], serial_in};
		   end else begin
		      temp_out <= {serial_in, temp_out[NUM_BITS-1:1]};
		   end
		end	
	end	
     end
  assign parallel_out = temp_out;

 endmodule
