// $Id: $
// File name:   bresenCircle.sv
// Created:     11/29/2016
// Author:      Vignesh Karthikeyan
// Lab Section: 337-07
// Version:     1.0  Initial Design Entry
// Description: bresenham's circle algorithm
