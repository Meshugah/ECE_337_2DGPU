//Module:
//Author(s): Noah Petersen
