//Module: Output Logic - This probably should be broken up more but oh well
//Authors